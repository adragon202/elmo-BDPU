module mean( a, b, mn);
	//input declaration
	input a, b;
	//output declaration
	output mn;
	//port data types
	wire a, b, mn;
	//code starts here

endmodule //addbit