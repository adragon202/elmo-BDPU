module squareroot( a, sqrt);
	//input declaration
	input a;
	//output declaration
	output sqrt;
	//port data types
	wire a, sqrt;
	//code starts here

endmodule //addbit