module product( a, b, prod);
	//input declaration
	input a, b;
	//output declaration
	output prod;
	//port data types
	wire a, b, prod;
	//code starts here

endmodule //addbit