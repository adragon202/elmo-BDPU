module square( a, sqr);
	//input declaration
	input a;
	//output declaration
	output sqr;
	//port data types
	wire a, sqr;
	//code starts here
	product P1(a(a),b(a),prod(sqr));

endmodule //addbit