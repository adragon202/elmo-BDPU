module bram( a, b, out);
	//input declaration
	input a, b;
	//output declaration
	output out;
	//port data types
	wire a, b, out;
	//code starts here

endmodule //addbit