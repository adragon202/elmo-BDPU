// main 	Top level of design, incorporating all other modules in some degree
//			This is where all components are connected and cores multiplied

//Libraries
module main();

endmodule //main