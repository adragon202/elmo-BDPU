module test;

	initial begin
		# 0 clk = 0;
		# 0 rst = 1;
		# 0 en = 0;
		//Sum of all zeroes
		// # 0 a[0] = 32'h0;
		// # 0 a[1] = 32'h0;
		// # 0 a[2] = 32'h0;
		// # 0 a[3] = 32'h0;
		// # 0 a[4] = 32'h0;
		// # 0 a[5] = 32'h0;
		// # 0 a[6] = 32'h0;
		// # 0 a[7] = 32'h0;
		// # 0 a[8] = 32'h0;
		// # 0 a[9] = 32'h0;
		// # 0 a[10] = 32'h0;
		// # 0 a[11] = 32'h0;
		// # 0 a[12] = 32'h0;
		// # 0 a[13] = 32'h0;
		// # 0 a[14] = 32'h0;
		// # 0 a[15] = 32'h0;
		// # 0 sum_expected = 32'h0;
		//Sum of max values
		// # 0 a[0] = 32'hffffffff;
		// # 0 a[1] = 32'hffffffff;
		// # 0 a[2] = 32'hffffffff;
		// # 0 a[3] = 32'hffffffff;
		// # 0 a[4] = 32'hffffffff;
		// # 0 a[5] = 32'hffffffff;
		// # 0 a[6] = 32'hffffffff;
		// # 0 a[7] = 32'hffffffff;
		// # 0 a[8] = 32'hffffffff;
		// # 0 a[9] = 32'hffffffff;
		// # 0 a[10] = 32'hffffffff;
		// # 0 a[11] = 32'hffffffff;
		// # 0 a[12] = 32'hffffffff;
		// # 0 a[13] = 32'hffffffff;
		// # 0 a[14] = 32'hffffffff;
		// # 0 a[15] = 32'hffffffff;
		// # 0 sum_expected = 32'hffffffff; //TODO: float Sums to 0x81ffffff
		//==================================
		//=============INT TESTS============
		//==================================
		// Sum of all 1's 00000001
		// # 0 a[0] = 32'h00000001;
		// # 0 a[1] = 32'h00000001;
		// # 0 a[2] = 32'h00000001;
		// # 0 a[3] = 32'h00000001;
		// # 0 a[4] = 32'h00000001;
		// # 0 a[5] = 32'h00000001;
		// # 0 a[6] = 32'h00000001;
		// # 0 a[7] = 32'h00000001;
		// # 0 a[8] = 32'h00000001;
		// # 0 a[9] = 32'h00000001;
		// # 0 a[10] = 32'h00000001;
		// # 0 a[11] = 32'h00000001;
		// # 0 a[12] = 32'h00000001;
		// # 0 a[13] = 32'h00000001;
		// # 0 a[14] = 32'h00000001;
		// # 0 a[15] = 32'h00000001;
		// # 0 sum_expected = 32'h00000010;
		//Sum to 1 from top
		// # 0 a[0] = 32'h00000001;
		// # 0 a[1] = 32'h0;
		// # 0 a[2] = 32'h0;
		// # 0 a[3] = 32'h0;
		// # 0 a[4] = 32'h0;
		// # 0 a[5] = 32'h0;
		// # 0 a[6] = 32'h0;
		// # 0 a[7] = 32'h0;
		// # 0 a[8] = 32'h0;
		// # 0 a[9] = 32'h0;
		// # 0 a[10] = 32'h0;
		// # 0 a[11] = 32'h0;
		// # 0 a[12] = 32'h0;
		// # 0 a[13] = 32'h0;
		// # 0 a[14] = 32'h0;
		// # 0 a[15] = 32'h0;
		// # 0 sum_expected = 32'h00000001;
		//Sum to 1 from bottom
		// # 0 a[0] = 32'h0;
		// # 0 a[1] = 32'h0;
		// # 0 a[2] = 32'h0;
		// # 0 a[3] = 32'h0;
		// # 0 a[4] = 32'h0;
		// # 0 a[5] = 32'h0;
		// # 0 a[6] = 32'h0;
		// # 0 a[7] = 32'h0;
		// # 0 a[8] = 32'h0;
		// # 0 a[9] = 32'h0;
		// # 0 a[10] = 32'h0;
		// # 0 a[11] = 32'h0;
		// # 0 a[12] = 32'h0;
		// # 0 a[13] = 32'h0;
		// # 0 a[14] = 32'h0;
		// # 0 a[15] = 32'h00000001;
		// # 0 sum_expected = 32'h00000001;
		//Sum a range of values
		// # 0 a[0] = 32'h33d6bf95; //869711765 +
		// # 0 a[1] = 32'h3f800000; //1065353216 +
		// # 0 a[2] = 32'h40000000; //1073741824 +
		// # 0 a[3] = 32'h40658106; //1080393990 +
		// # 0 a[4] = 32'h4080075f; //1082132319 +
		// # 0 a[5] = 32'h40ac6a7f; //1085041279 +
		// # 0 a[6] = 32'h40c00000; //1086324736 +
		// # 0 a[7] = 32'h40ff74bc; //1090483388 +
		// # 0 a[8] = 32'h44480000; //1145569280 +
		// # 0 a[9] = 32'h42b49a03; //1119132163 +
		// # 0 a[10] = 32'h41200000; //1092616192 +
		// # 0 a[11] = 32'h4133367a; //1093875322 +
		// # 0 a[12] = 32'h41463127; //1095119143 +
		// # 0 a[13] = 32'h41528f5c; //1095929692 +
		// # 0 a[14] = 32'h4808b800; //1208530944 +
		// # 0 a[15] = 32'h3c75c28f; //1014350479
		// # 0 sum_expected = 32'h070F32C4; //17298305732 (118436548)
		//Sum a range of negative values
		// # 0 a[0] = 32'hb3d6bf95; //-1277771883 +
		// # 0 a[1] = 32'hbf800000; //-1082130432 +
		// # 0 a[2] = 32'hc0000000; //-1073741824 +
		// # 0 a[3] = 32'hc0658106; //-1067089658 +
		// # 0 a[4] = 32'hc080075f; //-1065351329 +
		// # 0 a[5] = 32'hc0ac6a7f; //-1062442369 +
		// # 0 a[6] = 32'hc0c00000; //-1061158912 +
		// # 0 a[7] = 32'hc0ff74bc; //-1057000260 +
		// # 0 a[8] = 32'hc4480000; //-1001914368 +
		// # 0 a[9] = 32'hc2b49a03; //-1028351485 +
		// # 0 a[10] = 32'hc1200000; //-1054867456 +
		// # 0 a[11] = 32'hc133367a; //-1053608326 +
		// # 0 a[12] = 32'hc1463127; //-1052364505 +
		// # 0 a[13] = 32'hc1528f5c; //-1051553956 +
		// # 0 a[14] = 32'hc808b800; //-938952704 +
		// # 0 a[15] = 32'hbc75c28f; //-1133133169
		// # 0 sum_expected = 32'h78f0cd3c; //-17061432636 (overflow) (given (0x070f32c4)
		//Sum a mix of positive and negative values
		// # 0 a[0] = 32'hb3d6bf95; //-1277771883 +
		// # 0 a[1] = 32'h3f800000; //1065353216 +
		// # 0 a[2] = 32'hc0000000; //-1073741824 +
		// # 0 a[3] = 32'h40658106; //1080393990 +
		// # 0 a[4] = 32'hc080075f; //-1065351329 +
		// # 0 a[5] = 32'h40ac6a7f; //1085041279 +
		// # 0 a[6] = 32'hc0c00000; //-1061158912 +
		// # 0 a[7] = 32'h40ff74bc; //1090483388 +
		// # 0 a[8] = 32'hc4480000; //-1001914368 +
		// # 0 a[9] = 32'h42b49a03; //1119132163 +
		// # 0 a[10] = 32'hc1200000; //-1054867456 +
		// # 0 a[11] = 32'h4133367a; //1093875322 +
		// # 0 a[12] = 32'hc1463127; //-1052364505 +
		// # 0 a[13] = 32'h41528f5c; //1095929692 +
		// # 0 a[14] = 32'hc808b800; //-938952704 +
		// # 0 a[15] = 32'h3c75c28f; //1014350479
		// # 0 sum_expected = 32'h070F32C4; //118436548
		//==================================
		//============FLOAT TESTS===========
		//==================================
		//Sum of all 1's 3f800000
		# 0 a[0] = 32'h3f800000;
		# 0 a[1] = 32'h3f800000;
		# 0 a[2] = 32'h3f800000;
		# 0 a[3] = 32'h3f800000;
		# 0 a[4] = 32'h3f800000;
		# 0 a[5] = 32'h3f800000;
		# 0 a[6] = 32'h3f800000;
		# 0 a[7] = 32'h3f800000;
		# 0 a[8] = 32'h3f800000;
		# 0 a[9] = 32'h3f800000;
		# 0 a[10] = 32'h3f800000;
		# 0 a[11] = 32'h3f800000;
		# 0 a[12] = 32'h3f800000;
		# 0 a[13] = 32'h3f800000;
		# 0 a[14] = 32'h3f800000;
		# 0 a[15] = 32'h3f800000;
		# 0 sum_expected = 32'h41800000;
		//Sum to 1 from top
		// # 0 a[0] = 32'h3f800000;
		// # 0 a[1] = 32'h0;
		// # 0 a[2] = 32'h0;
		// # 0 a[3] = 32'h0;
		// # 0 a[4] = 32'h0;
		// # 0 a[5] = 32'h0;
		// # 0 a[6] = 32'h0;
		// # 0 a[7] = 32'h0;
		// # 0 a[8] = 32'h0;
		// # 0 a[9] = 32'h0;
		// # 0 a[10] = 32'h0;
		// # 0 a[11] = 32'h0;
		// # 0 a[12] = 32'h0;
		// # 0 a[13] = 32'h0;
		// # 0 a[14] = 32'h0;
		// # 0 a[15] = 32'h0;
		// # 0 sum_expected = 32'h3f800000;
		//Sum to 1 from bottom
		// # 0 a[0] = 32'h0;
		// # 0 a[1] = 32'h0;
		// # 0 a[2] = 32'h0;
		// # 0 a[3] = 32'h0;
		// # 0 a[4] = 32'h0;
		// # 0 a[5] = 32'h0;
		// # 0 a[6] = 32'h0;
		// # 0 a[7] = 32'h0;
		// # 0 a[8] = 32'h0;
		// # 0 a[9] = 32'h0;
		// # 0 a[10] = 32'h0;
		// # 0 a[11] = 32'h0;
		// # 0 a[12] = 32'h0;
		// # 0 a[13] = 32'h0;
		// # 0 a[14] = 32'h0;
		// # 0 a[15] = 32'h3f800000;
		// # 0 sum_expected = 32'h3f800000;
		//Sum a range of values
		// # 0 a[0] = 32'h33d6bf95; //0.0000001 +
		// # 0 a[1] = 32'h3f800000; //1 +
		// # 0 a[2] = 32'h40000000; //2 +
		// # 0 a[3] = 32'h40658106; //3.586 +
		// # 0 a[4] = 32'h4080075f; //4.0009 +
		// # 0 a[5] = 32'h40ac6a7f; //5.388000004 (5.388) +
		// # 0 a[6] = 32'h40c00000; //6 +
		// # 0 a[7] = 32'h40ff74bc; //7.983 +
		// # 0 a[8] = 32'h44480000; //800 +
		// # 0 a[9] = 32'h42b49a03; //90.3008007 +
		// # 0 a[10] = 32'h41200000; //10 +
		// # 0 a[11] = 32'h4133367a; //11.2008 +
		// # 0 a[12] = 32'h41463127; //12.387 +
		// # 0 a[13] = 32'h41528f5c; //13.16 +
		// # 0 a[14] = 32'h4808b800; //140000.00001 +
		// # 0 a[15] = 32'h3c75c28f; //0.015
		// # 0 sum_expected = 32'h4809a9c1; //140967.021511 (140967.02)
		//Sum a range of negative values
		// # 0 a[0] = 32'hb3d6bf95; //-0.0000001 +
		// # 0 a[1] = 32'hbf800000; //-1 +
		// # 0 a[2] = 32'hc0000000; //-2 +
		// # 0 a[3] = 32'hc0658106; //-3.586 +
		// # 0 a[4] = 32'hc080075f; //-4.0009 +
		// # 0 a[5] = 32'hc0ac6a7f; //-5.388000004 (5.388) +
		// # 0 a[6] = 32'hc0c00000; //-6 +
		// # 0 a[7] = 32'hc0ff74bc; //-7.983 +
		// # 0 a[8] = 32'hc4480000; //-800 +
		// # 0 a[9] = 32'hc2b49a03; //-90.3008007
		// # 0 a[10] = 32'hc1200000; //-10 +
		// # 0 a[11] = 32'hc133367a; //-11.2008 +
		// # 0 a[12] = 32'hc1463127; //-12.387 +
		// # 0 a[13] = 32'hc1528f5c; //-13.16 +
		// # 0 a[14] = 32'hc808b800; //-140000.00001 +
		// # 0 a[15] = 32'hbc75c28f; //-0.015
		// # 0 sum_expected = 32'hc809a9c1; //-140967.021511 (140967.02)
		//Sum a mix of positive and negative values
		// # 0 a[0] = 32'hb3d6bf95; //-0.0000001 +
		// # 0 a[1] = 32'h3f800000; //1 +
		// # 0 a[2] = 32'hc0000000; //-2 +
		// # 0 a[3] = 32'h40658106; //3.586 +
		// # 0 a[4] = 32'hc080075f; //-4.0009 +
		// # 0 a[5] = 32'h40ac6a7f; //5.388000004 (5.388) +
		// # 0 a[6] = 32'hc0c00000; //-6 +
		// # 0 a[7] = 32'h40ff74bc; //7.983 +
		// # 0 a[8] = 32'hc4480000; //-800 +
		// # 0 a[9] = 32'h42b49a03; //90.3008007
		// # 0 a[10] = 32'hc1200000; //-10 +
		// # 0 a[11] = 32'h4133367a; //11.2008 +
		// # 0 a[12] = 32'hc1463127; //-12.387 +
		// # 0 a[13] = 32'h41528f5c; //13.16 +
		// # 0 a[14] = 32'hc808b800; //-140000.00001 +
		// # 0 a[15] = 32'h3c75c28f; //0.015
		// # 0 sum_expected = 32'hc8096187; //-140678.111765 (-140678.11) (gave -140701.77)
		# 11 rst = 0;
		# 10 en = 1;
		# 300 $stop;
	end

	/* Pulse input */
	reg clk, rst, en;
	reg [31:0] a[0:15];
	reg [31:0] sum_expected;
	wire [31:0] sum;
	wire [31:0] in0, in1;
	wire [31:0] sums[0:3];
	wire rdy;

	always
		#5 clk  = !clk;

	accumulator #(.FLOAT(1)) accum_1(.EN(en), .clk(clk), .rst(rst),
		.vals({a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15]}), 
		.sum(sum), .rdy(rdy),
		.in0(in0), .in1(in1), .sum0(sums[0]), .sum1(sums[1]), .sum2(sums[2]), .sum3(sums[3]));

	initial
		$monitor("%g\t rst(%b), en(%b), SUM(a[0](0x%h)) = sum(?0x%h?)(0x%h) (%b) (in0(0x%h) + in1(0x%h) = sum0(0x%h), sum1(0x%h), sum2(0x%h), sum3(0x%h))",
				$time, rst, en, a[0], sum_expected, sum, rdy, in0, in1, sums[0], sums[1], sums[2], sums[3]);

endmodule //test