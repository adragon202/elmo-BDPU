-- main

architecture main of main is
begin
	core: 	WORK.sub-core generic map()
			port map();
	bram:	WORK.sub-bram generic map()
			port map();
	run: process
	begin

	end process;
end main;

